module Map (
    input rst,
    input clk,
    output reg [0:899] map //20*15 //(h+20*v)*3 (每格有3bit可使用)
);
    parameter NONE = 3'd0;
    parameter LINE = 3'd1;
    parameter TERMINAL = 3'd2;

    always @(posedge clk or posedge rst) begin
        if(rst) begin
            map <= { //最外圈須維持NONE
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0
            };
        end
        else map <= map; //之後做調整
    end
    
endmodule