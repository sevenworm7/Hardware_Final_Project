module Map (
    input rst,
    input clk,
    input [2:0] state,
    output reg [0:899] map //20*15 //(h+20*v)*3 (每格有3bit可使用)
);
    parameter NONE = 3'd0;
    parameter LINE = 3'd1;
    parameter TERMINAL = 3'd2;

    initial begin
        map <= {
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0
            };
    end

    always @(posedge clk or posedge rst) begin
        if(rst || state==3'b010) begin
            map <= { //最外圈須維持NONE
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd2, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0
            };
        end else if(state==3'b011) begin//win scene
            map <={
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0,
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0,
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0,
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0
            };
        end else if(state== 3'b100) begin
            map <={
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd0, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0,
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0,
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0,
                3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0
            };
        end
    end
    
endmodule