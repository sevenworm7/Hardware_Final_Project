module Led (
    input rst,
	input clk,
    input div_hsec,
    input state,
    input [2:0] curr_hp,
    output [15:0] LED
);
    
endmodule