module Seven_segment (
    input rst,
    input div_15,
    input [15:0] num,
    output [6:0] DISPLAY,
    output [3:0] DIGIT
);

    
endmodule