module Led (
    input rst,
	input clk,
    output [15:0] led
);
    
endmodule