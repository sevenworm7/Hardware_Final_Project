module Screen (
    input rst,
    input div_2,
    output [3:0] vgaRed,    
    output [3:0] vgaGreen,
    output [3:0] vgaBlue,   
    output hsync,           
    output vsync       
);
//參考 lab6 的範例2
    
endmodule