module Charactor (
    input rst,
    input clk,
    input key_num,
    input key,
    output charactor_posi
);
    
endmodule