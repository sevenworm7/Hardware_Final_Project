module Voice (
    input rst,
    input clk,
    input div_22,
    output audio_mclk, 
    output audio_lrck, 
    output audio_sck,  
    output audio_sdin 
);
//參考lab7
    
endmodule